----------------------------------------------------------------------
-- Created by Microsemi SmartDesign Sun Jun  7 23:40:11 2020
-- Parameters for CoreTimer
----------------------------------------------------------------------


LIBRARY ieee;
   USE ieee.std_logic_1164.all;
   USE ieee.std_logic_unsigned.all;
   USE ieee.numeric_std.all;

package coreparameters is
    constant FAMILY : integer := 19;
    constant INTACTIVEH : integer := 1;
    constant WIDTH : integer := 32;
end coreparameters;
